import "DPI-C" function void set_gpr_ptr(input longint regfile_0,input longint regfile_1,input longint regfile_2,input longint regfile_3,input longint regfile_4,input longint regfile_5,input longint regfile_6,input longint regfile_7,input longint regfile_8,input longint regfile_9,input longint regfile_10,input longint regfile_11,input longint regfile_12,input longint regfile_13,input longint regfile_14,input longint regfile_15,input longint regfile_16,input longint regfile_17,input longint regfile_18,input longint regfile_19,input longint regfile_20,input longint regfile_21,input longint regfile_22,input longint regfile_23,input longint regfile_24,input longint regfile_25,input longint regfile_26,input longint regfile_27,input longint regfile_28,input longint regfile_29,input longint regfile_30,input longint regfile_31);
module gpr_ptr(input clock,
	input reset,
	input [63:0] regfile_0,
       	input [63:0] regfile_1, 
	input [63:0] regfile_2,
	input [63:0] regfile_3,
	input [63:0] regfile_4,
	input [63:0] regfile_5,
	input [63:0] regfile_6,
	input [63:0] regfile_7,
	input [63:0] regfile_8,
	input [63:0] regfile_9,
	input [63:0] regfile_10,
	input [63:0] regfile_11,
	input [63:0] regfile_12,
	input [63:0] regfile_13,
	input [63:0] regfile_14,
	input [63:0] regfile_15,
	input [63:0] regfile_16,
	input [63:0] regfile_17,
	input [63:0] regfile_18,
	input [63:0] regfile_19,
	input [63:0] regfile_20,
	input [63:0] regfile_21,
	input [63:0] regfile_22,
	input [63:0] regfile_23,
	input [63:0] regfile_24,
	input [63:0] regfile_25,
	input [63:0] regfile_26,
	input [63:0] regfile_27,
	input [63:0] regfile_28,
	input [63:0] regfile_29,
	input [63:0] regfile_30,
	input [63:0] regfile_31
);

	always @(*)
		set_gpr_ptr(regfile_0, regfile_1, regfile_2, regfile_3, regfile_4,regfile_5,regfile_6,regfile_7,regfile_8,regfile_9,regfile_10,regfile_11,regfile_12,regfile_13,regfile_14,regfile_15,regfile_16,regfile_17,regfile_18,regfile_19,regfile_20,regfile_21,regfile_22,regfile_23,regfile_24,regfile_25,regfile_26,regfile_27,regfile_28,regfile_29,regfile_30,regfile_31);
endmodule
